`timescale 1ns/1ps

module and_gate_tb;

    reg a, b;
    wire y;

    and_gate dut (
        .a(a),
        .b(b),
        .y(y)
    );

    initial begin
        $display("A B | Y");
        a = 0; b = 0; #10;
        a = 0; b = 1; #10;
        a = 1; b = 0; #10;
        a = 1; b = 1; #10;
        $finish;
    end

    initial begin
        $monitor("%b %b | %b", a, b, y);
    end
    initial begin
    $dumpfile("and_gate.vcd");
    $dumpvars(0, and_gate_tb);
end


endmodule
